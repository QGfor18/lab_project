`timescale 1ns / 1ps

module top(
    input wire clk,             
    input wire uart_rx,         
    output wire uart_tx,        
    input wire [7:0] key,       // key[3:0] ��Ӧ SW3-SW0
    output wire [7:0] led,      // led[3:0] ��ʾ�洢״̬
    input wire uart_rx_rst_n,   // ��λ T5
    input wire btn_print_v1     // ��ӡ��ť V1
);
    
    // �ź�����
    wire [7:0] rx_data;
    wire rx_done;
    wire [7:0] tx_data;
    wire tx_start;
    wire tx_busy;
    
    // �����ź�
    wire btn_print_stable;
    
    // === ʵ���� ����ģ�� ===
    debounce u_db (
        .clk(clk),
        .rst_n(uart_rx_rst_n),
        .btn_in(btn_print_v1),
        .btn_out(btn_print_stable)
    );
    
    // UART RX
    uart_rx #( .CLK_FREQ(100_000_000), .BAUD_RATE(115200) ) u_rx (
        .clk(clk), .rst_n(uart_rx_rst_n),
        .rx(uart_rx), .rx_data(rx_data), .rx_done(rx_done)
    );
    
    // UART TX
    uart_tx #( .CLK_FREQ(100_000_000), .BAUD_RATE(115200) ) u_tx (
        .clk(clk), .rst_n(uart_rx_rst_n),
        .tx_start(tx_start), .tx_data(tx_data),
        .tx(uart_tx), .tx_busy(tx_busy)
    );
    
    // === ���Ŀ���ģ�� ===
    matrix_io_ctrl u_ctrl (
        .clk(clk), .rst_n(uart_rx_rst_n),
        .rx_data(rx_data), .rx_done(rx_done),
        .tx_data(tx_data), .tx_start(tx_start), .tx_busy(tx_busy),
        
        // �ؼ������޸�
        .print_trigger(btn_print_stable), // ʹ��������� V1 �ź�
        .sw_select(key[3:0]),             // ʹ�� SW0-SW3 ѡ���������
        .led(led[3:0])                    // LED0-3 ��ʾ�洢״̬
    );
    
    // δʹ�õ� LED Ϩ��
    assign led[7:4] = 4'b0000;
    
endmodule
`timescale 1ns / 1ps

module debounce(
    input wire clk,       // 100MHz
    input wire rst_n,
    input wire btn_in,    // ԭʼ��������
    output reg btn_out    // ������İ������
);

    // 20ms ����ʱ��: 100MHz * 0.02s = 2,000,000
    parameter CNT_MAX = 2_000_000;
    
    reg [20:0] cnt;
    reg btn_d1, btn_d2;
    
    // ��ʱ��������ģ���������̬
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            btn_d1 <= 0;
            btn_d2 <= 0;
        end else begin
            btn_d1 <= btn_in;
            btn_d2 <= btn_d1;
        end
    end

    // �����������߼�
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            cnt <= 0;
            btn_out <= 0;
        end else begin
            // �������״̬�仯�����ü�����
            if(btn_d2 != btn_out) begin
                cnt <= cnt + 1;
                if(cnt >= CNT_MAX) begin
                    btn_out <= btn_d2; // ״̬�ȶ����������
                    cnt <= 0;
                end
            end else begin
                cnt <= 0; // ״̬δ�䣬����
            end
        end
    end
endmodule